/****************************
        >Title:async_fifo

****************************/
module async_fifo();

